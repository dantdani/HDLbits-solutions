module top_module ( input x, input y, output z );
    // simple xnor gate!
    xnor simple(z, x, y);
​
endmodule
