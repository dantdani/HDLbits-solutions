module top_module (
    input in,
    output out);
