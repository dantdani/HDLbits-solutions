module top_module (input x, input y, output z);

endmodule

module A (input x, input y, output z);

endmodule

module B (input x, input y, output z);

endmodule
