module top_module ( 
    input [15:0] a, b,
    input cin,
    output cout,
    output [15:0] sum );

endmodule
