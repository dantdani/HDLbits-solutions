module top_module( 
    input a, b, sel,
    output out ); 

endmodule
