module top_module ( input x, input y, output z );
