module top_module( 
    input [399:0] a, b,
    input cin,
    output cout,
    output [399:0] sum );
