module top_module (input x, input y, output z);
    wire o1, o2, o3, o4;
    
    A ia1 (x, y, o1);
    B ib1 (x, y, o2);
    A ia2 (x, y, o3);
    B ib2 (x, y, o4);
    
    assign z = (o1 | o2) ^ (o3 & o4);
endmodule

module A (input x, input y, output z);
    assign z = (x^y) & x;
endmodule

module B (input x, input y, output z);
    assign z = ~(x^y);
endmodule
