module top_module (
    output out);
