module top_module (
    input in1,
    input in2,
    output out);
    nor mu_nor(out, in1,in2);
​
endmodule
