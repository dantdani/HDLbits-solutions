module top_module( 
    input a, b, cin,
    output cout, sum );

endmodule
