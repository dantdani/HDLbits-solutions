module top_module( 
    input [2:0] in,
    output [1:0] out );

endmodule
